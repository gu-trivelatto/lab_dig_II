--------------------------------------------------------------------
-- Arquivo   : interface_hcsr04_tb.vhd
-- Projeto   : Experiencia 4 - Interface com sensor de distancia
--------------------------------------------------------------------
-- Descricao : testbench para circuito de interface com HC-SR04 
--
--             1) array de casos de teste contém valores de  
--                largura de pulso de echo do sensor
-- 
--------------------------------------------------------------------
-- Revisoes  :
--     Data        Versao  Autor             Descricao
--     19/09/2021  1.0     Edson Midorikawa  versao inicial
--------------------------------------------------------------------
--
library ieee;
use ieee.std_logic_1164.all;

entity interface_hcsr04_tb is
end entity;

architecture tb of interface_hcsr04_tb is
  
  -- Componente a ser testado (Device Under Test -- DUT)
  component interface_hcsr04
    port (
            clock, reset:    in  std_logic;
            medir:           in  std_logic;
            echo:            in  std_logic;
            trigger:         out std_logic;
            medida:          out std_logic_vector(11 downto 0);
            pronto:          out std_logic;
            db_estado:       out std_logic_vector(3 downto 0);
            db_dist0:        out std_logic_vector (6 downto 0);
            db_dist1:        out std_logic_vector (6 downto 0);
            db_dist2:        out std_logic_vector (6 downto 0);
            db_medir:        out std_logic; 
            db_reset:        out std_logic;
            db_trigger:      out std_logic; 
            db_echo:         out std_logic;
            db_estado_sseg : out std_logic_vector (6 downto 0)
    );
  end component;
  
  -- Declaração de sinais para conectar o componente a ser testado (DUT)
  --   valores iniciais para fins de simulacao (GHDL ou ModelSim)
  signal clock_in:            std_logic := '0';
  signal reset_in:            std_logic := '0';
  signal medir_in:            std_logic := '0';
  signal echo_in:             std_logic := '0';
  signal medida_out:          std_logic_vector (11 downto 0) := x"000";
  signal trigger_out:         std_logic := '0';
  signal pronto_out:          std_logic := '0';
  signal db_estado_out:       std_logic_vector (3 downto 0) := "0000";
  signal db_dist0_out :       std_logic_vector (6 downto 0) := "0000000";
  signal db_dist1_out :       std_logic_vector (6 downto 0) := "0000000";
  signal db_dist2_out :       std_logic_vector (6 downto 0) := "0000000";
  signal db_medir_out :       std_logic := '0';
  signal db_reset_out :       std_logic := '0';
  signal db_trigger_out :     std_logic := '0';
  signal db_echo_out :        std_logic := '0';
  signal db_estado_sseg_out : std_logic_vector (6 downto 0) := "0000000";

  -- Configurações do clock
  signal keep_simulating: std_logic := '0'; -- delimita o tempo de geração do clock
  constant clockPeriod:   time := 20 ns;    -- clock de 50MHz
  
  -- Array de casos de teste
  type caso_teste_type is record
      id    : natural; 
      tempo : integer;     
  end record;

  type casos_teste_array is array (natural range <>) of caso_teste_type;
  constant casos_teste : casos_teste_array :=
      (
        (1, 5882),  -- 5882us (100cm)
        (2, 4353)   -- 4353us (74cm)
        -- inserir aqui outros casos de teste (inserir "," na linha anterior)
      );

  signal larguraPulso: time := 1 ns;

begin
  -- Gerador de clock: executa enquanto 'keep_simulating = 1', com o período
  -- especificado. Quando keep_simulating=0, clock é interrompido, bem como a 
  -- simulação de eventos
  clock_in <= (not clock_in) and keep_simulating after clockPeriod/2;
  
  -- Conecta DUT (Device Under Test)
  dut: interface_hcsr04
       port map( clock=>      clock_in,
                 reset=>      reset_in,
                 medir=>      medir_in,
                 echo=>       echo_in,
                 trigger=>    trigger_out,
                 medida=>     medida_out,
                 pronto=>     pronto_out,
                 db_estado => db_estado_out,
                 db_dist0 => db_dist0_out,
                 db_dist1 => db_dist1_out,
                 db_dist2 => db_dist2_out,
                 db_medir => db_medir_out,
                 db_reset => db_reset_out,
                 db_trigger => db_trigger_out,
                 db_echo => db_echo_out,
                 db_estado_sseg => db_estado_sseg_out
      );

  -- geracao dos sinais de entrada (estimulos)
  stimulus: process is
  begin
  
    assert false report "Inicio das simulacoes" severity note;
    keep_simulating <= '1';
    
    ---- valores iniciais ----------------
    medir_in <= '0';
    echo_in  <= '0';

    ---- inicio: reset ----------------
    wait for 2*clockPeriod;
    reset_in <= '1'; 
    wait for 2 us;
    reset_in <= '0';
    wait until falling_edge(clock_in);

    ---- espera de 100us
    wait for 100 us;

    ---- loop pelos casos de teste
    for i in casos_teste'range loop
        -- 1) determina largura do pulso echo
        assert false report "Caso de teste " & integer'image(casos_teste(i).id) & ": " &
            integer'image(casos_teste(i).tempo) & "us" severity note;
        larguraPulso <= casos_teste(i).tempo * 1 us; -- caso de teste "i"

        -- 2) envia pulso medir
        wait until falling_edge(clock_in);
        medir_in <= '1';
        wait for 5*clockPeriod;
        medir_in <= '0';
     
        -- 3) espera por 400us (tempo entre trigger e echo)
        wait for 400 us;
     
        -- 4) gera pulso de echo (largura = larguraPulso)
        echo_in <= '1';
        wait for larguraPulso;
        echo_in <= '0';
     
        -- 5) espera final da medida
      	wait until pronto_out = '1';
        assert false report "Fim do caso " & integer'image(casos_teste(i).id) severity note;
     
        -- 6) espera entre casos de tese
        wait for 100 us;

    end loop;

    ---- final dos casos de teste da simulacao
    assert false report "Fim das simulacoes" severity note;
    keep_simulating <= '0';
    
    wait; -- fim da simulação: aguarda indefinidamente (não retirar esta linha)
  end process;

end architecture;
